library verilog;
use verilog.vl_types.all;
entity Memory is
    port(
        I_CLOCK         : in     vl_logic;
        I_LOCK          : in     vl_logic;
        I_Opcode        : in     vl_logic_vector(7 downto 0);
        I_PC            : in     vl_logic_vector(15 downto 0);
        I_IR            : in     vl_logic_vector(31 downto 0);
        I_R15PC         : in     vl_logic_vector(15 downto 0);
        I_DestRegIdx    : in     vl_logic_vector(3 downto 0);
        I_DestVRegIdx   : in     vl_logic_vector(5 downto 0);
        I_DestValue     : in     vl_logic_vector(15 downto 0);
        I_CCValue       : in     vl_logic_vector(2 downto 0);
        I_VecSrc1Value  : in     vl_logic_vector(63 downto 0);
        I_VecDestValue  : in     vl_logic_vector(63 downto 0);
        I_EX_Valid      : in     vl_logic;
        I_MARValue      : in     vl_logic_vector(15 downto 0);
        I_MDRValue      : in     vl_logic_vector(15 downto 0);
        I_RegWEn        : in     vl_logic;
        I_VRegWEn       : in     vl_logic;
        I_CCWEn         : in     vl_logic;
        I_GPUStallSignal: in     vl_logic;
        O_LOCK          : out    vl_logic;
        O_Opcode        : out    vl_logic_vector(7 downto 0);
        O_IR            : out    vl_logic_vector(31 downto 0);
        O_PC            : out    vl_logic_vector(15 downto 0);
        O_R15PC         : out    vl_logic_vector(15 downto 0);
        O_DestRegIdx    : out    vl_logic_vector(3 downto 0);
        O_DestVRegIdx   : out    vl_logic_vector(5 downto 0);
        O_LEDR          : out    vl_logic_vector(9 downto 0);
        O_LEDG          : out    vl_logic_vector(7 downto 0);
        O_HEX0          : out    vl_logic_vector(6 downto 0);
        O_HEX1          : out    vl_logic_vector(6 downto 0);
        O_HEX2          : out    vl_logic_vector(6 downto 0);
        O_HEX3          : out    vl_logic_vector(6 downto 0);
        O_CCValue       : out    vl_logic_vector(2 downto 0);
        O_VecSrc1Value  : out    vl_logic_vector(63 downto 0);
        O_VecDestValue  : out    vl_logic_vector(63 downto 0);
        O_DestValue     : out    vl_logic_vector(15 downto 0);
        O_MEM_Valid     : out    vl_logic;
        O_RegWEn        : out    vl_logic;
        O_VRegWEn       : out    vl_logic;
        O_CCWEn         : out    vl_logic
    );
end Memory;
