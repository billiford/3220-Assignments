library verilog;
use verilog.vl_types.all;
entity Decode is
    port(
        I_CLOCK         : in     vl_logic;
        I_LOCK          : in     vl_logic;
        I_PC            : in     vl_logic_vector(15 downto 0);
        I_IR            : in     vl_logic_vector(31 downto 0);
        I_FE_Valid      : in     vl_logic;
        I_WriteBackRegIdx: in     vl_logic_vector(3 downto 0);
        I_WriteBackVRegIdx: in     vl_logic_vector(5 downto 0);
        I_WriteBackData : in     vl_logic_vector(15 downto 0);
        I_CCValue       : in     vl_logic_vector(2 downto 0);
        I_WriteBackPC   : in     vl_logic_vector(15 downto 0);
        I_WriteBackPCEn : in     vl_logic;
        I_VecSrc1Value  : in     vl_logic_vector(63 downto 0);
        I_VecSrc2Value  : in     vl_logic_vector(63 downto 0);
        I_VecDestValue  : in     vl_logic_vector(63 downto 0);
        I_RegWEn        : in     vl_logic;
        I_VRegWEn       : in     vl_logic;
        I_CCWEn         : in     vl_logic;
        I_EDDestRegIdx  : in     vl_logic_vector(3 downto 0);
        I_EDDestVRegIdx : in     vl_logic_vector(5 downto 0);
        I_EDDestWrite   : in     vl_logic;
        I_EDDestVWrite  : in     vl_logic;
        I_MDDestRegIdx  : in     vl_logic_vector(3 downto 0);
        I_MDDestVRegIdx : in     vl_logic_vector(5 downto 0);
        I_MDDestWrite   : in     vl_logic;
        I_MDDestVWrite  : in     vl_logic;
        I_EDCCWEn       : in     vl_logic;
        I_MDCCWEn       : in     vl_logic;
        I_GPUStallSignal: in     vl_logic;
        O_LOCK          : out    vl_logic;
        O_PC            : out    vl_logic_vector(15 downto 0);
        O_Opcode        : out    vl_logic_vector(7 downto 0);
        O_IR            : out    vl_logic_vector(31 downto 0);
        O_Src1Value     : out    vl_logic_vector(15 downto 0);
        O_Src2Value     : out    vl_logic_vector(15 downto 0);
        O_DestRegIdx    : out    vl_logic_vector(3 downto 0);
        O_DestVRegIdx   : out    vl_logic_vector(5 downto 0);
        O_Idx           : out    vl_logic_vector(1 downto 0);
        O_Imm           : out    vl_logic_vector(15 downto 0);
        O_DepStallSignal: out    vl_logic;
        O_BranchStallSignal: out    vl_logic;
        O_CCValue       : out    vl_logic_vector(2 downto 0);
        O_VecSrc1Value  : out    vl_logic_vector(63 downto 0);
        O_VecSrc2Value  : out    vl_logic_vector(63 downto 0);
        O_DE_Valid      : out    vl_logic
    );
end Decode;
